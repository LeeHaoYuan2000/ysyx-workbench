module DIV(
    input [63:0] src1,
    input [63:0] src2,
    input control,   //0 is src1 / src2 , 1 is src1 % src2
    output [63:0] result_out
    );

assign
endmodule