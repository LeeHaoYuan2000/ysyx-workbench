module CSR(
    input [31:0] Instr,
    
);
endmodule
