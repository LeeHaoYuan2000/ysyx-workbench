module SEXT(
    input [31:0] Instr,
    input [] ControlUnit,
    output [63:0] sext
);

endmodule
